netcdf initial_from_climatology {                           
dimensions:                                                 
	time = UNLIMITED ;                                         
	s_rho = 50 ;                                               
	eta_rho = 441 ;                                            
	xi_rho = 204 ;                                             
	eta_u = 441 ;                                              
	xi_u = 203 ;                                               
	eta_v = 440 ;                                              
	xi_v = 204 ;                                               
variables:                                                  
	double time(time) ;                                        
		time:long_name = "HYCOM climatology time" ;               
		time:units = "seconds since 2003-12-31 00:00:00" ;        
		time:calendar = "gregorian" ;                             
		time:field = "time, scalar, series" ;                     
	double ocean_time(time) ;                                  
		ocean_time:long_name = "HYCOM climatology time" ;         
		ocean_time:units ="seconds since 2003-12-31 00:00:00" ;   
		ocean_time:calendar = "gregorian" ;                       
		ocean_time:field = "time, scalar, series" ;               
	float temp(time, s_rho, eta_rho, xi_rho) ;                 
		temp:long_name = "potential temperature" ;                
		temp:units = "Celsius" ;                                  
		temp:time = "time" ;                                      
		temp:field = "temp, scalar, series" ;                     
	float salt(time, s_rho, eta_rho, xi_rho) ;                 
		salt:long_name = "salinity" ;                             
		salt:units = "PSU" ;                                      
		salt:time = "time" ;                                      
		salt:field = "salt, scalar, series" ;                     
	float u(time, s_rho, eta_u, xi_u) ;                        
		u:long_name = "u-velocity component" ;                    
		u:units = "meter second-1" ;                              
		u:time = "time" ;                                         
		u:field = "u, scalar, series" ;                           
	float ubar(time, eta_u, xi_u) ;                            
		ubar:long_name = "ubar-velocity component" ;              
		ubar:units = "meter second-1" ;                           
		ubar:time = "time" ;                                      
		ubar:field = "ubar, scalar, series" ;                     
	float v(time, s_rho, eta_v, xi_v) ;                        
		v:long_name = "v-velocity component" ;                    
		v:units = "meter second-1" ;                              
		v:time = "time" ;                                         
		v:field = "v, scalar, series" ;                           
	float vbar(time, eta_v, xi_v) ;                            
		vbar:long_name = "vbar-velocity component" ;              
		vbar:units = "meter second-1" ;                           
		vbar:time = "time" ;                                      
		vbar:field = "vbar, scalar, series" ;                     
	float zeta(time, eta_rho, xi_rho) ;                        
		zeta:long_name = "sea surface height" ;                   
		zeta:units = "meter" ;                                    
		zeta:time = "time" ;                                      
		zeta:field = "zeta, scalar, series" ;                     
                                                            
// global attributes:                                       
		:type = "ROMS initial condition file" ;                   
		:history = "Generated with initial_from_climatology.f90 " ;         
		:title ="ROMS ini file for the domain /scratch/rw408/Input_COAWST/Ang5km_V2/Angola_grid_5km_V2.nc" ;                       
		:source = "HYCOM" ;                                       
		:source_url = "Inputs from HYCOM files: /scratch/cdenamie/HYCOM/CONGO" ;                          
}                                                           
