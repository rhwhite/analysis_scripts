netcdf climatology_file {                                   
dimensions:                                                 
	time = UNLIMITED ;                                         
	s_rho = 35 ;                                               
	eta_rho = 463 ;                                            
	xi_rho = 305 ;                                             
	eta_u = 463 ;                                              
	xi_u = 304 ;                                               
	eta_v = 462 ;                                              
	xi_v = 305 ;                                               
variables:                                                  
	float salt(time, s_rho, eta_rho, xi_rho) ;                 
		salt:long_name = "salinity" ;                             
		salt:units = "PSU" ;                                      
		salt:time = "time" ;                                      
		salt:field = "salt, scalar, series" ;                     
	float temp(time, s_rho, eta_rho, xi_rho) ;                 
		temp:long_name = "potential temperature" ;                
		temp:units = "Celsius" ;                                  
		temp:time = "time" ;                                      
		temp:field = "temp, scalar, series" ;                     
	double time(time) ;                                        
		time:long_name = "HYCOM climatology time" ;               
		time:units = "seconds since 2003-12-31 00:00:00" ;        
		time:calendar = "gregorian" ;                             
		time:field = "time, scalar, series" ;                     
	float u(time, s_rho, eta_u, xi_u) ;                        
		u:long_name = "u-velocity component" ;                    
		u:units = "meter second-1" ;                              
		u:time = "time" ;                                         
		u:field = "u, scalar, series" ;                           
	float ubar(time, eta_u, xi_u) ;                            
		ubar:long_name = "ubar-velocity component" ;              
		ubar:units = "meter second-1" ;                           
		ubar:time = "time" ;                                      
		ubar:field = "ubar, scalar, series" ;                     
	float v(time, s_rho, eta_v, xi_v) ;                        
		v:long_name = "v-velocity component" ;                    
		v:units = "meter second-1" ;                              
		v:time = "time" ;                                         
		v:field = "v, scalar, series" ;                           
	float vbar(time, eta_v, xi_v) ;                            
		vbar:long_name = "vbar-velocity component" ;              
		vbar:units = "meter second-1" ;                           
		vbar:time = "time" ;                                      
		vbar:field = "vbar, scalar, series" ;                     
	float zeta(time, eta_rho, xi_rho) ;                        
		zeta:long_name = "sea surface height" ;                   
		zeta:units = "meter" ;                                    
		zeta:time = "time" ;                                      
		zeta:field = "zeta, scalar, series" ;                     
                                                            
// global attributes:                                       
		:type = "ROMS climatology file" ;                         
		:title ="ROMS Climatology file generated for the domain /scratch/rw408/Input_COAWST/Nam5km_V1/Namibia_grid_5km_V1.nc" ;                             
		:source = "HYCOM" ;                                       
		:source_url = "Inputs from HYCOM files: /scratch/cdenamie/HYCOM/CONGO." ;                         
}                                                           
